----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:40:46 02/23/2017 
-- Design Name: 
-- Module Name:    ROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
--use IEEE.STD_LOGIC_ARITH.all;
use IEEE.NUMERIC_STD.all;

entity ROM is
    Port ( clk : 				in  STD_LOGIC;
           mem_address : 	in  STD_LOGIC_VECTOR (15 downto 0);
           data : 			out  STD_LOGIC_VECTOR (15 downto 0));
end ROM;

architecture Behavioral of ROM is

    type ROM_TYPE is array (0 to 41) of std_logic_vector (7 downto 0);

    constant rom_content : ROM_TYPE := (
	 
	 -- FINAL TEST 1 -- 0 to 41
	"00100100","00000011", -- LOADIMM.lower 3
	"00100111","10111000", -- MOV 	R6, R7
	"00100100","00000001", -- LOADIMM.lower 1
	"00100111","01111000", -- MOV 	R5, R7
	"01000010","00000000", -- IN 		R0
	"00000010","01000110", -- ADD 	R1, R0 + R6
	"00000110","10000000", -- MUL 	R2, R0 * R0
	"00000110","11001001", -- MUL 	R3, R1 * R1
	"00000100","11011010", -- SUB 	R3, R3 - R2
	"00100011","01011000", -- STORE 	M[R5], R3
	"00000010","10000001", -- ADD 	R2, R0, R1
	"00100011","00010000", -- STORE 	M[R4], R2
	"00100000","10100000", -- LOAD 	R2, M[R4]
	"00100000","11101000", -- LOAD 	R3, M[R5]
	"00000100","11011010", -- SUB 	R3, R3 - R2	 
	"00001110","11000000", -- TEST 	R3
	"10000100","00000010", -- BRRZ	2
	"00000101","10110101", -- SUB 	R6, R6 - R5
	"10000111","01000100", -- BR 		R5, 4
	"01000000","10000000", -- OUT 	R2
	"10000001","11101011"); -- BRR	-21	

		-- FINAL TEST 2 -- 0 to 27
--	"00100100","00000001", -- LOADIMM.lower 1
--	"00100111","01111000", -- MOV 	R5, R7
--	"00100110","01101000", -- MOV 	R1, R5
--	"00100111","10101000", -- MOV 	R6, R5
--	"00001011","10000001", -- SHL 	R6, 1
--	"01000010","00000000", -- IN 		R0
--	"00000110","01001000", -- MUL 	R1, R1 * R0
--	"00000100","00000101", -- SUB 	R0, R0 - R5
--	"00000101","00000110", -- SUB 	R4, R0 - R6 
--	"00001111","00000000", -- TEST 	R4
--	"10000010","00000001", -- BRRN	1
--	"10000111","10000100", -- BR 		R6, 4
--	"01000000","01000000", -- OUT 	R1
--	"10000001","11110010"); -- BRR	-14	
		
	 
	 
	 -- FORMAT B TEST 2 --
--	"01000010","00000000", -- IN R0 , 02  -- This example tests the branching capabilities of the design.No data dependencies.
--	"01000010","01000000", -- IN R1 , 03  -- The values to be loaded into the corresponding resgister.
--	"01000010","10000000", -- IN R2 , 01
--	"01000010","11000000", -- IN R3 , 05  --  End of initialization
--	"01000011","00000000", -- IN R4 , 00
--	"01000011","01000000", -- IN R5 , 01  -- for absolute branching
--	"01000011","10000000", -- IN R6 , 05  -- r6 is counter for the loop and indicates the number of times the loop is done.
--	"01000011","11000000", -- IN R7 , 00
--	"10001101","00000001", -- BR.SUB R4, 1 -- Go to the subroutine
--	"10000001","11111111", -- BRR -1     -- Infinite loop (the end of the program)
--	"00000010","10001101", -- ADD R2, R1, R5  -- Start of the subroutine. It runs for 5 times. R2 <-- R1 + 1
--	"00000101","10110101", -- SUB R6, R6, R5  -- R6 <-- R6 - 1   The counter for the loop.
--	"00001111","10000000", -- TEST R6         -- Set the z flag for the branch decision
--	"10001011","00000001", -- BR.z R4, 1      -- If r6 is zero, jump out of the loop. 
--	"10000001","11111011", -- BRR -5		-- If not jump to the start of the subroutine.	 
--	"10001110","00000000", -- RET
--	"00000000","00000000"); -- NOP	 
	
--	"01000010","00000000",
--	"00000000","00000000",
--	"00000000","00000000",
--	"00000000","00000000",
--	"00000000","00000000",
--	"00000000","00000000",
--	"00000000","00000000",
--	"00000000","00000000",
--	"01000000","00000000",
--	"00000000","00000000",
--	"00000000","00000000",
--	"00000000","00000000",
--	"00000000","00000000",
--	"00000000","00000000",
--	"00000000","00000000",
--	"00000000","00000000",
--	"00000000","00000000"); -- NOP	
	 
	 -- FORMAT L TEST --
--	"00100100","00001111", -- LOADIMM.LOWER #15
--	"00100101","00000101", -- LOADIMM.UPPER #5
--	"00100110","01111000", -- MOV R1, R7
--	"00100100","00000110", -- LOADIMM.LOWER #6
--	"00100101","00000000", -- LOADIMM.UPPER #0
--	"00100110","10111000", -- MOV R2, R7
--	"00100010","10001000", -- STORE R2, R1
--	"00100000","11010000", -- LOAD R3, R1
--	"00000000","00000000", -- NOP
--	"00000000","00000000", -- NOP
--	"00000000","00000000"); -- NOP
	 
--		"01000010",
--		"01000000",  -- IN r1
--		"01000010",
--		"10000000",  -- IN r2
--		"01000010",
--		"11000000",  -- IN r3	
--		"00000100",
--		"11001010",  -- SUB r3, r1, r2
--		"00001010",
--		"10000010",  -- SHL r3, 2
--		"00000110",
--		"10001011",  -- MUL r2, r1, r3
--		"00001110",
--		"11000000",	 -- TEST r3
--		"10000011",
--		"11111100",	 -- BRN -4 
--		"00000010",
--		"11001010",  -- ADD r3, r1, r2
--		"00000000",
--		"00000000",	 -- NOP
--		"00000000",
--		"00000000"); -- NOP	
		
		-- Test Branching BRN, BRZ - Use r1 = 1, r2 = 2, r3 = 5 --
--		"01000010",
--		"01000000",  -- IN r1
--		"01000010",
--		"10000000",  -- IN r2
--		"01000010",
--		"11000000",  -- IN r3	
--		"00000100",
--		"10001011",  -- SUB r2, r1, r3
--		"00000010",
--		"10010001",  -- ADD r2, r2, r1
--		"00001110",
--		"10000000",	 -- TEST r2
--		"10001000",
--		"01111101",	 -- BRN r1 -3 
--		"00001110",
--		"10000000",	 -- TEST r2
--		"10001010",
--		"01111011",	 -- BRZ r1 -5
--		"00000000",
--		"00000000",	 -- NOP
--		"00000000",
--		"00000000"); -- NOP	
		
		-- Test Branching BRSUB, Return --
--		"01000010",
--		"01000000",  -- IN r1
--		"00000000",
--		"00000000",	 -- NOP
--		"10001100",
--		"01000011",	 -- BRSUB r1 +3 	
--		"00000010",
--		"01001001",  -- ADD r1, r1, r1
--		"00000000",
--		"00000000",	 -- NOP	
--		"00000000",
--		"00000000",  -- NOP	
--		"00000000",
--		"00000000",	 -- NOP	
--		"00000000",
--		"00000000",	 -- NOP	
--		"00000000",
--		"00000000",	 -- NOP
--		"10001110",
--		"00000000",	 -- RET	
--		"00000000",
--		"00000000"); -- NOP	
		
		-- Test Memory --
--		"01000010",
--		"01000000",  -- IN r1
--		"01000010",
--		"10000000",  -- IN r2
--		"00100010",
--		"01010000",	 -- STORE r2 > M[r1] 	
--		"00100001",
--		"10001000",	 -- LOAD M[r1] > r6
--		"00100010",
--		"10110000",	 -- STORE r6 > M[r2]		
--		"00000000",
--		"00000000",	 -- NOP 		
--		"00000000",
--		"00000000",	 -- NOP			
--		"00000000",
--		"00000000",	 -- NOP	
--		"00000000",
--		"00000000",	 -- NOP
--		"00000000",
--		"00000000",	 -- NOP	
--		"00000000",
--		"00000000"); -- NOP	
		
begin

	data <= rom_content(to_integer(unsigned(mem_address))) & rom_content(to_integer(unsigned(mem_address))+ 1);

end Behavioral;

